library IEEE;
use ieee.std_logic_1164.all;


ENTITY dec_7seg IS
   PORT(W : IN std_logic_vector(3 downto 0);
		F : OUT std_logic_vector(5 downto 0));       	
END dec_7seg;

architecture behavior OF dec_7seg IS
begin
end behavior;